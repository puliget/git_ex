fb.log
